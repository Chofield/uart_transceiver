%TSD-Header-###%9l3����3� 2H  �           @  ����.   �P �v*�	)XN��-�뇞����4��QK�!h*��qE���<�9S��!!��!�����V�hfaI��Pt>U�3ث9(�7pa)XN��-�뇞�M��4��P��!h섦q����,�9R��!1���!����V���XI)XNQ��뇶�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        {	�úi���J���b���.��xؙ��-,��J����+��I'W��B��IL��w=��I���c��?̸����s�[�[\�����v�~xk���=6e�����JQLS�A���?�Ult��=���4�hoׄ}��В�0[	�{�R�Is24��k�RQ�Q6/��8���7ܱABR��1ϼ�(x�v���«�yB#O�T��쐀2��5f�ƈ�5�kՄ�wü�Z]�'0���.*�^T�� :��y�EZ<����m��E�&�5�8ϼʛ��A�Ʊ�.�m�3;��A���؞<22GL2�(b����N�I;������Z���k?`T�KU��Î��@>ۊ0�.�ȺM�`\RC�y����ƺV~���tjf&O��|�$201rj���\��s��Pyd�& #� �� RR0��0�V�M"y=Dj���:��ff<J�K�����;5e��>o.�$ȸ�pޠ�n����9�b�ɹ`̇��3^e�0����ѯ���o�@�
8�O�����'�U��'qt�V�a������9��&�1�ܸ������Ų�o�۹�f�Ò���W�I5���#�T����CE�����m������7Ī%��s�[��ԼDQ���U����դR �(���;��o�i��(h���1KX�H�.]��IcqY��!�[����L�j���t0��l[J�4�,���u�1x��E��&�C�~�2zw�_y`���������C���X0�[���C�cSݨ�%�X=F0�8V���-��#���@���Lx�
�k�c����1��bH�X�^^v�8͍OG��y�/op����n��uVX욗R�Ɛ��MJR����e����VTmco�Q�[�7���� ٞo��o�v�=A'�8d�:�^5�J�(�����5��|���s�جO|[�b����X��iO��,
)���T8�y8%�ZӉ�x���kT��%����X�U�_�!���D$�[���jrT����4�bԜ\�.�c�@Q2�/ɼoc�q�Gfh�u_�\YUr�ɩ��7��_��#�,���g2mj�O�:� Z`�������R� ApW�Zi��	[B�+��g�/I ��r	u_X�DЫMX��	S��\@�ͅ,�~����޲�6�:f3��!��{<o�z�\��2k3̠�����Z�Y�%�4�6�����a ��1U�d%��CӇ��3̵�<jtr�,P�b`��
P�'��ڶ��A�7o�� pp_w$̿�l%��8���|N��bW���"���i�߿��g�t�'�E�+]*�����\�!���A���t�"�n_A�12�z�E�FK�j�SM���x���'\/>+Tc��%�㇔QP7��[���/��9���b��TxM� �5��n��]�5�6�� ��lı�Wn;�7�VƳj"��!���㩘7�q6�<z��ꙡ�?���T	g�ŏ��=��{�����û?��������<�'�w�V���@M���5�̪|���+n~�%M��o:J6%;��g"�LQ�F�ȍ��PU�N��`C7�i%��i���8]�V��.��+sҟ��W�h������)n)�2�x���m*����S�����S]���w%t`Y �k#J3�~�9�>�@�D;Xֲ��{{l�~�պD�u\��=�>�q�	�r�~�'\��V���f(:��TB3�оa�#F�Q��b4h��c���zE9�}���Q���w}4�f���\,�����V��UD��ٟ����gFa��;\0����������"�i�5d��֤u�Mrm�aJP*�y�'g��Z�5�p76xQ�0[2pghe�A
�M��<PG`�c^Ĳ;A��-�����{��({��ȅj�W`G}m���j�[�y�[tΞ�Mf��+�M�y���,��{�|=O��s��I��/@#�T�.ыM�&�Ɣ���T�tM�����W[�mkw��bh��%n���U�����$,d�9��_�):~2Vs����v�f#ڶ�2}@��7�s� ���}���v=GH�BR2�$�B�x~���eϐfwv���j��]�n�\��K��ٚ�e���:׀��Y�4wȹ��.�	>>.��7��\�8̎ߤ�Y&�յ�ϋ�5@%���D�xt(}N<�8m����=��M�^ЦZ��-�׉]��3U�sY ~������3�"�+����6IU���W�Lq���̼vN�e�b��M��]
� (��9h.NcJ�	�x�q�m V����)�ȐBI��ֿ�5���{�(�4�Q;�A���Bק���8�
śS�5<�#��[qIq�c�8Uh�aN�	���։'+w!E1F7���'�0]�Y��C]?������Wj��R>�d��Q=o��9�?C̰��o�v,�oI��vyL��7��!���P�T�+����,YA�{ۥ���o9j�����"T��}?�s4W�_cX�舮����Y��Z7:KX?�ՙ�PJ/8bbU �S��f�+�Hv�!�:WmE���{M޽����!����r�z���Z�����0�t����;�R���*P%O�X��:n>�&���w/C���I�s����쌎�d�'�:��O/,����n�5;����ݢ��A !��tF�kN�J��ă�t�|�Z'U���<(+���/�+@;⫙S������ᚿ;q� Y�*\= BW\g^{��C�O���{7���s��.�y%��MĄlvm�d=~%4�> ��[�;��x��d(�������
�$��>���_</jOu�=�����
j!�LODC��.���S�B�����p\�����D&�S���߆�  4q���Y�N֯-��+毐�H���}�u1��85�Ƅ����H*m�dp*L�����'�]/o
 ��geXcM[��D�Z��`���z��d/̥�F~��C�V�uØ��wq���=-؋T=>iLо��)�T�T�u`�H\�\(�aM��
,�$w�o�#\8F]�9O�ָq��E��h_�%��X�@ưp��nEE���ُ����(r�3���K��@������j�G(NG��C�~�5c"��:
�i���lt�avU �I\��D�|�G��⚹�g��`�۩>t&�Z�5y��ޱ�0�ج,�q�u낔��v��BL��p%����ġE=���캠Zq�k]�!�K+������pij����ڞ�>�Z�����К��^��S�s7�H�İ�<��F����n�����t;���Z�}P�[Sꑒ���$u�MA�&��ps�AbQ"~��/���ƚ\���P�49yn�L6�,�Av�`#�=#�ni-#�_B����v�8I�*5+0�_�$��R����_e+�Ⱦ R�?�gү���?�7�o;Z���	�c�H�0#㇬aEU�Jh����;M�q�$Bc�X�uv�m�E)x}��R�#+����.��hn_?ydud��%�1����d������e��|�R�Ŏ9�9W���h,���b7E������"��E�rN���&Ϲ�|g�)�VbS�帿g8�A޼��2�KQ�k:��ƞ�o�&�j���6��9ƅ�X��ń|V�7g�c�}�	���g):~��w�3V�|��&�a@��	���,��s��P��C�R{�v4�n���6g"�|X �h�l�ڮL��eW��=�T(����R��U{<��i ���{��R׆5�
쬹�������$?��>�wѺ,\S�P�1����N[��؉�nR��>�ӹp)��3s%y�<�J/^O�����=AQ]�o���[������j?��cc�M4t�3
��I�w_���v���0mY�6��/�Wk3�hS/뇊��.�W���4��c'�Lne���߾	�"��rCg��i+�V��ٺ̬�\��s'���&,bڠ@��[3�9Q�H���$��v��*�f���a�r��� �L�Zp�`���t�
EUfz����e��w�L;���